LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY deco7Seg IS 
PORT(
numero : IN INTEGER RANGE 0 TO 9;
HEX : OUT STD_LOGIC_VECTOR (7 DOWNTO 0) 
);
END deco7seg;
ARCHITECTURE prueba OF deco7seg IS 
BEGIN
	WITH numero SELECT
		HEX<= "11000000" WHEN 0,
				"11111001" WHEN 1,
				"10100100" WHEN 2,
				"10110000" WHEN 3,
				"10011001" WHEN 4,
				"10010010" WHEN 5,
				"10000010" WHEN 6,
				"11111000" WHEN 7,
				"10000000" WHEN 8,
				"10010000" WHEN 9,
				"11111111" WHEN OTHERS;


END prueba;